
`define DELAY 20
module ALUtb();
	reg [31:0] a, b;
    reg [3:0] ALUControl;
    wire zeroes;

    wire [31:0] result;
	
alu potaot (result,zeroes,a,b,ALUControl)	;
initial begin
// AND tests, start
    ALUControl = 3'b000;
	a = 32'b00000000000000000000000000000000;
    b = 32'b00000000000000000000000000000000;
#`DELAY;
    a = 32'b11111111111111111111111111111111;
    b = 32'b11111111111111111111111111111111;
#`DELAY;
    a = 32'b00000000000000000000000000001100;
    b = 32'b00000000000000000000000000001010;
#`DELAY;
// AND tests, end.

// OR tests, start
    ALUControl = 3'b001;
	a = 32'b00000000000000000000000000000000;
    b = 32'b00000000000000000000000000000000;
#`DELAY;
    a = 32'b11111111111111111111111111111111;
    b = 32'b11111111111111111111111111111111;
#`DELAY;
    a = 32'b00000000000000000000000000001100;
    b = 32'b00000000000000000000000000001010;
#`DELAY;
// OR tests, end.

// ADD tests, start
    ALUControl = 3'b010;
	a = 32'b00000000000000000000000000000000;
    b = 32'b00000000000000000000000000000000;
#`DELAY;
    a = 32'b00000000000000000000000000001100;
    b = 32'b00000000000000000000000000001010;
#`DELAY;
// ADD tests, end.

// SUBSTRACT tests, start
    ALUControl = 3'b110;
	a = 32'b11111111111111111111111111111111;
    b = 32'b11111111111111111111111111111111;
#`DELAY;
    a = 32'b00000000000000000000000000001100;
    b = 32'b00000000000000000000000000001010;
#`DELAY;
    a = 32'b00000000000000000000000000001010;
    b = 32'b00000000000000000000000000001100;
#`DELAY;
// SUBSTRACT tests, end.

// XOR tests, start
    ALUControl = 3'b011;
	a = 32'b00000000000000000000000000000000;
    b = 32'b00000000000000000000000000000000;
#`DELAY;
    a = 32'b11111111111111111111111111111111;
    b = 32'b11111111111111111111111111111111;
#`DELAY;
    a = 32'b00000000000000000000000000001100;
    b = 32'b00000000000000000000000000001010;
#`DELAY;
// XOR tests, end.

end

initial begin
	$monitor("a=%32b, b=%32b, ALUControl=%3b, result=%32b, zero=%1b",a, b, ALUControl, result, zeroes);
end

endmodule